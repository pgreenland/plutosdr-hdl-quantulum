`timescale 1ns / 1ps

module util_upack2_timestamp_tb;
    reg clk;
    reg reset;
    wire reset_upack;
    reg [63:0] timestamp;
    reg [31:0] timestamp_every;
    reg s_axis_valid;
    wire s_axis_ready;
    reg s_axis_xfer_req;
    reg [63:0] s_axis_data;
    wire m_axis_valid;
    wire m_axis_ready;
    wire [63:0] m_axis_data;

    util_upack2_timestamp #( 
        .NUM_OF_CHANNELS (4),
        .SAMPLE_DATA_WIDTH (16),
        .SAMPLES_PER_CHANNEL (1)
    ) uut (
        .dma_clk(clk),
        .dac_clk(clk),
        .reset(reset),
        .reset_upack(reset_upack),
        .timestamp(timestamp),
        .timestamp_every(timestamp_every),
        .s_axis_valid(s_axis_valid),
        .s_axis_ready(s_axis_ready),
        .s_axis_xfer_req(s_axis_xfer_req),
        .s_axis_data(s_axis_data),
        .m_axis_valid(m_axis_valid),
        .m_axis_ready(m_axis_ready),
        .m_axis_data(m_axis_data)
    );

    always begin
        // Toggle clock
        #1 clk = ~clk;
    end

    always @(posedge clk) begin
        // Increment timestamp
        timestamp <= timestamp + 1;
    end 

    // Test mode
    localparam MODE_READ_VECTORS = 0;
    localparam MODE_WRITE_VECTORS = 1;
    reg mode = MODE_READ_VECTORS;

    // Test vector - unpack reset + data bits
    reg [64:0] expected_outputs [0:35];

    integer i, j;
    reg ts_req;

    initial begin
        // Load test vectors
        if (mode == MODE_READ_VECTORS)
            $readmemb("util_upack2_timestamp_tv_vectors.mem", expected_outputs);

        // Reset signals
        clk = 'b0;
        reset = 'b1;
        timestamp = 'h0;
        timestamp_every = 'h0;
        s_axis_valid = 'b0;
        s_axis_xfer_req = 'b0;
        s_axis_data = 'h0;

        // De-assert reset
        @(posedge clk)
        reset <= 1'b0;

        // Wait for FIFO to come out of reset
        #164;

        // Reset sample counter
        j = 0;

        // Perform test with timestamping disabled, enabled and late, enabled and on time, enabled and early
        for (i = 0; i < 4; i = i + 1) begin
            // Set mode
            if (i == 0) begin
                // Timestamping disabled
                timestamp_every = 'h0;
            end else begin
                // Timestamping enabled
                timestamp_every = 'h4;
            end

            // Assert transfer request
            @(posedge clk)
            s_axis_xfer_req <= 'b1;

            // Iterate through test values
            ts_req = 'b1;
            while (j < ((i + 1) * 48)) begin          
                // Provide data on first step, or if ready asserted
                @(posedge clk)
                if (!s_axis_valid || s_axis_ready) begin
                    // Insert timestamp every x blocks
                    if (timestamp_every != 0 && ((j / 4) % timestamp_every == 0) && ts_req) begin
                        // Provide timestamp
                        case (i)
                            // Timestamp late
                            1: s_axis_data[63:0] <= timestamp;
                            // Timestamp on time
                            2: s_axis_data[63:0] <= timestamp + 1;
                            // Timestamp early
                            3: s_axis_data[63:0] <= timestamp + 2;
                        endcase

                        // Assert data valid
                        s_axis_valid <= 'b1;
                        
                        // Clear timestamp required
                        ts_req <= 'b0;
                    end else begin
                        // Provide record
                        s_axis_data[48+:16] <= j+4;
                        s_axis_data[32+:16] <= j+3;
                        s_axis_data[16+:16] <= j+2;
                        s_axis_data[0+:16] <= j+1;
                        s_axis_valid <= 'b1;
                
                        // Increment index
                        j = j + 4;

                        // Set timestamp required
                        ts_req <= 'b1;
                    end
                end
            end
           
            // Wait for final value to be consumed
            @(posedge clk)
            while (!s_axis_ready) begin
                #2;       
            end

            // Clear valid flag, reset data and deassert transfer request
            s_axis_data <= 'h0;
            s_axis_valid <= 'b0;
            s_axis_xfer_req <= 'b0;
            
            // Delay for clock cycle
            #2;
        end

        // Wait for reads to complete
        #32;

        // Write captured expected vectors out to file
        if (mode == MODE_WRITE_VECTORS)
            $writememb("util_upack2_timestamp_tv_vectors.mem", expected_outputs);

        // Got this far without error, all must be good
        $display("Test PASSED");

        // All done
        $finish;
    end
   
    // Wait for valid signal and print data
    integer expected_index = 0;
    always @(posedge clk) begin
        if (reset_upack) begin
            $display("Output: Reset");
        end

        if (m_axis_valid) begin
            // Dump data
            $display("Output: %h", m_axis_data);
        end

        if (reset_upack || m_axis_valid) begin
            // Compare to expected (or update expected)
            if (mode == MODE_READ_VECTORS) begin
                // Compare output to expected
                if (expected_outputs[expected_index] != {reset_upack, m_axis_valid ? m_axis_data : 64'h0}) begin
                    $error("Test FAILED, Expected: %b,%h got %b,%h",
                           expected_outputs[expected_index][64],
                           expected_outputs[expected_index][63:0],
                           reset_upack,
                           m_axis_valid ? m_axis_data : 64'h0);
                    $finish;
                end
            end else begin
                // Store output as expected         
                expected_outputs[expected_index] = {reset_upack, m_axis_valid ? m_axis_data : 64'h0};
            end          

            // Increment index
            expected_index = expected_index + 1;
        end
    end

    // For test purposes we'll accept data whenever we can get it
    assign m_axis_ready = m_axis_valid;
endmodule
